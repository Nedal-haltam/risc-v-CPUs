
`include "defs.h"

module HW_Interface(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,
	output		     [7:0]		HEX2,
	output		     [7:0]		HEX3,
	output		     [7:0]		HEX4,
	output		     [7:0]		HEX5,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// Arduino //////////
	inout 		    [15:0]		ARDUINO_IO,
	inout 		          		ARDUINO_RESET_N
);
`define CLK_BIT 15
reg [24:0] ClockDivider;
always@(posedge ADC_CLK_10) begin
	ClockDivider <= ClockDivider + 1'b1;
end
wire clk;
`define BUFFER_LEN 1025
reg [7:0] databuff [0 : `BUFFER_LEN - 1];

reg [31:0] index;
reg [7:0] DataOut;
reg done;

wire rst;
wire fillbuf;
wire datatrigger;

`define STR_LEN 10
integer i;
always@(posedge clk, posedge fillbuf) begin
	if (fillbuf) begin
		for (i = 0; i < `STR_LEN - 2; i = i + 1) begin : FillData
			databuff[i] = "a" + i;
		end
		databuff[`STR_LEN - 2] = "\n";
		databuff[`STR_LEN - 1] = 0;
	end
end

always@(posedge clk, posedge rst) begin
	if (rst) begin
		index = 0;
		DataOut = 0;
		done = 0;
	end
	else if (!done) begin
		done = (index >= `BUFFER_LEN) || (databuff[index] == 0);
		DataOut = databuff[index];
		index = index + 1'b1;
	end
end

assign datatrigger = (!done) ? rst | ~clk : 1'b0;
assign ARDUINO_IO[7:0] = DataOut;
assign ARDUINO_IO[8] = datatrigger;
assign ARDUINO_RESET_N = 1'b1;

assign clk = ClockDivider[`CLK_BIT];
assign rst = ~KEY[0];
assign fillbuf = ~KEY[1];

wire `BIT_WIDTH AddressBus, DataBusIn, DataBusOut;
wire [2:0] ControlBus;

CPU cpu_dut
(
	.InputClk(clk), 
	.rst(rst),
	.AddressBus(AddressBus),
	.DataBusIn(DataBusIn),
	.DataBusOut(DataBusOut),
	.ControlBus(ControlBus),
	.CyclesConsumed()
);

DataMemory MemoryModule
(
	.clock(~clk), 
    .MemReadEn(ControlBus[1]), 
    .MemWriteEn(ControlBus[2]),
	.AddressBus(AddressBus),
	.DataMemoryInput(DataBusOut),
	.DataMemoryOutput(DataBusIn)
);


endmodule

