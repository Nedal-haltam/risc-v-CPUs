
`include "defs.h"

module HW_Interface(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,
	output		     [7:0]		HEX2,
	output		     [7:0]		HEX3,
	output		     [7:0]		HEX4,
	output		     [7:0]		HEX5,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// Arduino //////////
	inout 		    [15:0]		ARDUINO_IO,
	inout 		          		ARDUINO_RESET_N
);

reg [24:0] ClockDivider;
always@(posedge ADC_CLK_10) begin
	ClockDivider <= ClockDivider + 1'b1;
end

reg `BIT_WIDTH offset;
reg [7:0] DataOut;
reg done;

wire clk;
wire rst;

wire exit_ecall;
wire write_ecall_finished;
wire write_ecall;
wire `BIT_WIDTH write_ecall_fd;
wire `BIT_WIDTH write_ecall_address;
wire `BIT_WIDTH write_ecall_len;
wire datatrigger;

wire `BIT_WIDTH AddressBus1, DataBusIn1, DataBusOut1, DataBusOut2, AddressBus2;
wire [10:0] ControlBus;
wire `BIT_WIDTH CyclesConsumed;

// FSM states
localparam IDLE    = 4'd0;
localparam SENDING = 4'd1;

reg [3:0] state;
always @(negedge clk or posedge rst) begin
    if (rst) begin
		done    <= 1'b1;
        offset  <= 0;
        DataOut <= 0;
        state   <= IDLE;
    end
	else begin
        case (state)

        IDLE: begin
			if (write_ecall) begin
				done    <= 1'b0;
				offset  <= 0;
				DataOut <= 0;
                state <= SENDING;
            end
			else begin
				done    <= 1'b1;
				offset  <= 0;
				DataOut <= 0;
				state <= IDLE;
			end
        end

        SENDING: begin
            if (offset < write_ecall_len) begin
				done <= 0;
                offset  <= offset + 1'b1;
                DataOut <= DataBusOut2[7:0];
            end
			else begin
				done <= 1'b1;
                offset  <= 0;
                DataOut <= 0;
				state <= IDLE;
            end
        end
        endcase
    end
end

CPU cpu_dut
(
	.InputClk(clk),
	.cpu_clk(cpu_clk),
	.rst(rst),
	.AddressBus(AddressBus1),
	.DataBusIn(DataBusIn1),
	.DataBusOut(DataBusOut1),
	.ControlBus(ControlBus),
	.CyclesConsumed(CyclesConsumed),

	.exit_ecall(exit_ecall),
	.write_ecall_finished(write_ecall_finished),
	.write_ecall(write_ecall),
	.write_ecall_fd(write_ecall_fd), // TODO: we should handle it, for now it is ignored
	.write_ecall_address(write_ecall_address),
	.write_ecall_len(write_ecall_len)
);

// TODO: use real altera dual-port ram 2 read / 2 write
DataMemory MemoryModule
(
	.rst(rst),
	.clock1(~clk),
	.loadtype1(ControlBus[6:3]),
	.storetype1(ControlBus[10:7]),
    .MemReadEn1(ControlBus[1]),
    .MemWriteEn1(ControlBus[2]),
	.AddressBus1(AddressBus1),
	.DataMemoryInput1(DataBusOut1),
	.DataMemoryOutput1(DataBusIn1),

	.clock2(clk),
	.loadtype2(`LOAD_BYTE), // TODO: drive the loadtype2, for now always byte
    .MemReadEn2(write_ecall),
    .MemWriteEn2(1'b0),
	.AddressBus2(write_ecall_address + offset),
	.DataMemoryInput2(),
	.DataMemoryOutput2(DataBusOut2)
);

assign datatrigger = (!done) ? (rst | clk) : (1'b0);
assign ARDUINO_IO[7:0] = DataOut;
assign ARDUINO_IO[8] = datatrigger;
assign ARDUINO_RESET_N = 1'b1;

assign write_ecall_finished = done;

assign clk = ClockDivider[17];
assign rst = ~KEY[0];

assign LEDR[0] = clk;
assign LEDR[1] = cpu_clk;
assign LEDR[2] = rst;
assign LEDR[3] = datatrigger;
assign LEDR[4] = done;
assign LEDR[5] = write_ecall_finished;
assign LEDR[6] = write_ecall;
assign LEDR[7] = exit_ecall;


endmodule

